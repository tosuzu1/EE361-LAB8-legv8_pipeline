// EE 361
// LEGLite 
// 
// The control module for LEGLite
//   The control will input the opcode value (3 bits)
//   then determine what the control signals should be
//   in the datapath
//  
//---------------------------------------------------------------
module Control(
     output logic reg2loc,
     output logic uncondbranch,
     output logic branch,
     output logic memread,
     output logic memtoreg,
     output logic [2:0] alu_select,
     output logic memwrite,
     output logic alusrc,
     output logic regwrite,
     input logic [3:0] opcode
     );


always_comb
	case(opcode)
	0:	// ADD
		begin
		reg2loc = 0;		//Pick 1st reg field
		uncondbranch = 0;	//Disable unconditional Branch
		branch = 0;   		//Disable Branch
		memread = 0;  		//Disable memory
		memtoreg = 0;		//Have ALU write to reg
		alu_select = 0; 	//Have ALU do an ADD
		memwrite = 0; 		//Disable memory
		alusrc = 0; 		//Read from register
		regwrite = 1;		//Write result to register
		end
	1:	// SUB
		begin
		reg2loc = 0;		//Pick 1st reg field
		uncondbranch = 0;	//Disable unconditional Branch
		branch = 0;   		//Disable Branch
		memread = 0;  		//Disable memory
		memtoreg = 0;		//Have ALU write to reg
		alu_select = 1; 	//Have ALU do an SUB
		memwrite = 0; 		//Disable memory
		alusrc = 0; 		//Read from register
		regwrite = 1;		//Write result to register
		end
	4:	// Branch
		begin
		reg2loc = 1;		//Pick 2nd reg field(Don't care for Branch)
		uncondbranch = 1;	//Enable unconditional Branch
		branch = 1;   		//Enable Branch
		memread = 0;  		//Disable memory
		memtoreg = 0;		//Have ALU write to reg
		alu_select = 0; 	//Have ALU do an ADD
		memwrite = 0; 		//Enable memory
		alusrc = 0; 		//Read from instruction
		regwrite = 0;		//Disable write to register
		end
	5:	// Load
		begin
		reg2loc = 1;		//Pick 2nd reg field(don't care for LDUR)
		uncondbranch = 0;	//Disable unconditional Branch
		branch = 0;   		//Disable Branch
		memread = 1;  		//Disable memory
		memtoreg = 1;		//Have Memory write to register
		alu_select = 0; 	//Have ALU do an ADD
		memwrite = 0; 		//Disable memory
		alusrc = 1; 		//Read from instruction
		regwrite = 1;		//Write result to register
		end
	6:	// Store
		begin
		reg2loc = 1;		//Pick 2nd reg field
		uncondbranch = 0;	//Disable unconditional Branch
		branch = 0;   		//Disable Branch
		memread = 0;  		//Disable memory
		memtoreg = 0;		//Have ALU write to reg
		alu_select = 0; 	//Have ALU do an ADD
		memwrite = 1; 		//Enable memory
		alusrc = 1; 		//Read from instruction
		regwrite = 0;		//Disable write to register
		end
	7:	// CBZ
		begin
		reg2loc = 1;		//Pick 2nd reg field
		uncondbranch = 0;	//Disable unconditional Branch
		branch = 1;   		//Enable Branch
		memread = 0;  		//Disable memory
		memtoreg = 0;		//Have ALU write to reg
		alu_select = 2; 	//Have ALU Cmp value to zero
		memwrite = 1; 		//Enable memory
		alusrc = 1; 		//Read from instruction
		regwrite = 0;		//Disable write to register
		end
	8:	// ADDI
		begin
		reg2loc = 0;		//Pick 2nd reg field
		uncondbranch = 0;	//Disable unconditional Branch
		branch = 0;   		//Disable Branch
		memread = 0;  		//Disable memory
		memtoreg = 0;		//Have ALU write to reg
		alu_select = 0; 	//Have ALU ADD
		memwrite = 0; 		//Enable memory
		alusrc = 1; 		//Read from instruction
		regwrite = 1;		//Disable write to register
		end
	9:	// ANDI
		begin
		reg2loc = 0;		//Pick 2nd reg field
		uncondbranch = 0;	//Disable unconditional Branch
		branch = 0;   		//Disable Branch
		memread = 0;  		//Disable memory
		memtoreg = 0;		//Have ALU write to reg
		alu_select = 4; 	//Have ALU ADD
		memwrite = 0; 		//Enable memory
		alusrc = 1; 		//Read from instruction
		regwrite = 1;		//Disable write to register
		end
	10:	// SUBI
		begin
		reg2loc = 0;		//Pick 2nd reg field
		uncondbranch = 0;	//Disable unconditional Branch
		branch = 0;   		//Disable Branch
		memread = 0;  		//Disable memory
		memtoreg = 0;		//Have ALU write to reg
		alu_select = 1; 	//Have ALU ADD
		memwrite = 0; 		//Enable memory
		alusrc = 1; 		//Read from instruction
		regwrite = 1;		//Disable write to register
		end
	default:
		begin
		reg2loc = 0;
		uncondbranch = 0;
		branch = 0;   
		memread = 0;   
		memtoreg = 0;  
		alu_select = 0; 
		memwrite = 0; 
		alusrc = 0;    
		regwrite = 0;
		end
	endcase

endmodule




